`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:36:36 11/17/2018 
// Design Name: 
// Module Name:    annh 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module annh(out,input1,input2);
input input1,input2;
output out;
wire input1,input2,out;
and And(out,input1,input2);
endmodule
